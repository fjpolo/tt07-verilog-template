/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_fjpolo_nes_apu (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // // All output pins must be assigned. If not used, assign to 0.
  // assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  // assign uio_out = 0;
  // assign uio_oe  = 0;

  simple_nes_apu my_apu(
    .simple_nes_apu_ui_in(ui_in),
    .simple_nes_apu_uo_out(uo_out),
    .simple_nes_apu_uio_in(uio_in),
    .simple_nes_apu_uio_out(uio_out),
    .simple_nes_apu_uio_oe(uio_oe),
    .simple_nes_apu_ena(ena),
    .simple_nes_apu_clk(clk),
    .simple_nes_apu_rst_n(rst_n)
  );

endmodule
